`include "defines.v"

module mem_control(
    input wire clk,
    input wire rst,
    input wire branch_interception,

    // interation with ram
    input wire[7:0] din_ram,
    output reg[7:0] dout_ram,
    output reg[`InstAddrBus] addr_ram,
    output reg wr_ram,
    
    output reg almost_available,
    output reg[`InstBus] inst,

    // interaction with if
    input wire[`InstAddrBus] inst_addr_i,
    output reg available,
    output reg[`InstAddrBus] inst_addr_o,

    // interaction with mem
    input wire datawr_i,
    input wire[`MemAddrBus] data_addr_i,
    input wire[`MemDataBus] data_i,
    input wire[1:0] data_cnf_i

);

    reg[2:0] cnt;
    reg[`InstAddrBus] addr;
    reg busy_inst;
    reg busy_mem;

    always @ (posedge clk) begin
        if (rst == `RstEnable) begin
            cnt <= 3'b110; //Since I begin with 0 here, the first instruction will step twice.
            almost_available <= `False;
            available <= `False;
            addr <= 0;
            dout_ram <= 0;
            wr_ram <= 0;
            inst <= 0;
            inst_addr_o <= 0;
            
        end else begin
            if (branch_interception) begin
                almost_available <= 1;
                cnt <= 0;
            end else if (cnt == 3'b000) begin
                case (data_cnf_i)
                2'b00: begin
                    addr <= inst_addr_i;
                    addr_ram <= inst_addr_i;
                    wr_ram <= 0;
                    almost_available <= `False;
                    available <= `False;
                    cnt <= cnt + 1;
                end
                2'b01: begin
                    addr <= data_addr_i;
                    addr_ram <= data_addr_i + 3;
                    dout_ram <= data_i;
                    wr_ram <= datawr_i;
                    almost_available <= `False;
                    available <= `False;
                    cnt <= cnt + 4;
                end
                2'b10: begin
                    addr <= data_addr_i;
                    addr_ram <= data_addr_i + 2;
                    dout_ram <= data_i;
                    wr_ram <= datawr_i;
                    almost_available <= `False;
                    available <= `False;
                    cnt <= cnt + 3;
                end
                2'b11: begin
                    addr <= data_addr_i;
                    addr_ram <= data_addr_i;
                    dout_ram <= data_i;
                    wr_ram <= datawr_i;
                    almost_available <= `False;
                    available <= `False;
                    cnt <= cnt + 1;
                end
                endcase
            end else if (cnt == 3'b001) begin
                addr_ram = addr + 1;
                cnt <= cnt + 1;
            end else if (cnt == 3'b010) begin
                inst[31:24] <= din_ram;
                addr_ram = addr + 2;
                cnt <= cnt + 1;
            end else if (cnt == 3'b011) begin
                inst[23:16] <= din_ram;
                addr_ram <= addr + 3;
                cnt <= cnt + 1;
            end else if (cnt == 3'b100) begin
                inst[15:8] <= din_ram;
                cnt <= cnt + 1;
            end else if (cnt == 3'b101) begin
                inst[7:0] <= din_ram;
                inst_addr_o <= addr;
                cnt <= 0;
                almost_available <= 1;
                available <= 1;
            end else if (cnt == 3'b110) begin
                almost_available <= 1;
                cnt <= 0;
            end

            /*
            if (cnt == 2'b00) begin
                inst[7:0] <= din_ram;
                addr_ram <= addr + 1;
                available <= `True;
                cnt <= 2'b01;
            end else if (cnt == 2'b01) begin
                inst[31:24] <= din_ram;
                addr_ram = addr + 2;
                available = `False;
                cnt <= 2'b10;
            end else if (cnt == 2'b10) begin
                inst[23:16] <= din_ram;
                addr_ram <= addr + 3;
                almost_available <= `True;
                cnt <= 2'b11;
            end else if (cnt == 2'b11) begin
                inst[15:8] <= din_ram;
                inst_addr_o <= addr; // Give back to PC
                almost_available <= `False;
                
                addr = inst_addr_i;
                addr_ram = addr;
                cnt = 2'b00;
                wr_ram = `Read;
            end
            */
        end
    end

endmodule